`timescale 1ns/10ps
`celldefine
module sg13g2_and2_2 (X, A, B);
	output X;
	input A, B;
	and (X, A, B);
endmodule
`endcelldefine
